module adcClock();
    

endmodule
