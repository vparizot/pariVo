module hardware_test(input  logic clk,
           input  logic [31:0] eqVals,
		   output logic ledTest);
		   
		   
	always_ff @(posedge clk)
		begin
			if (eqVals == 32'h12345678) ledTest <= 1;
			else ledTest <= 0;
				
		end
		
		
endmodule
